module sink (valid_ready_if.sink in);
  always_comb in.ready = 1'b1;
endmodule
