// Code your design here
`include "valid_ready_if.sv"
`include "diff.sv"
`include "sink.sv"
