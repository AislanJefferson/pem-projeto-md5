package diff_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "valid_ready_source_tx.svh"
  `include "valid_ready_source_driver.svh"
  `include "valid_ready_source_monitor.svh"
  `include "valid_ready_source_agent.svh"
  `include "valid_ready_source_seq_lib.svh"
  `include "valid_ready_sink_tx.svh"
  `include "valid_ready_sink_driver.svh"
  `include "valid_ready_sink_monitor.svh"
  `include "valid_ready_sink_agent.svh"
  `include "valid_ready_sink_seq_lib.svh"
  `include "bvm_comparator.svh"
  `include "diff_refmod.svh"

  `include "diff_env.svh"
  `include "diff_test.svh"
  `include "diff_sink_test.svh"
endpackage

