// Code your testbench here
// or browse Examples
`include "diff_pkg.sv"
`include "tb_diff.sv"
